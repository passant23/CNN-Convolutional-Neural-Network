`timescale 1ns / 1ps
module testbench_softmaxLayer();
reg clock;
reg reset;
parameter datawidth=32;
reg [datawidth-1:0] inputlayer [9:0][1][1]; 
wire [datawidth-1:0] outputlayer [9:0][1][1];


softmaxLayer S_Layer (clock,
reset,
inputlayer,
outputlayer
    );

initial begin
clock=1'b1;
reset=1'b0;
//0
inputlayer[0][0][0]=32'b00000000000000000000000000000000;
//1
inputlayer[1][0][0]=32'b00111111100000000000000000000000;
//-1
inputlayer[2][0][0]=32'b10111111100000000000000000000000;
//0.5
inputlayer[3][0][0]=32'b00111111000000000000000000000000;
//1
inputlayer[4][0][0]=32'b00111111100000000000000000000000;
//0.2
inputlayer[5][0][0]=32'b00111110010011001100110011001101;
//-0.5
inputlayer[6][0][0]=32'b10111111000000000000000000000000;
//0.3
inputlayer[7][0][0]=32'b00111110100110011001100110011010;
//0
inputlayer[8][0][0]=32'b00000000000000000000000000000000;
//0.7
inputlayer[9][0][0]=32'b00111111001100110011001100110011;
#600
//-1
inputlayer[0][0][0]=32'b10111111100000000000000000000000;
//0
inputlayer[1][0][0]=32'b00000000000000000000000000000000;
//-0.5
inputlayer[2][0][0]=32'b10111111000000000000000000000000;
//0.5
inputlayer[3][0][0]=32'b00111111000000000000000000000000;
//-0.66
inputlayer[4][0][0]=32'b10111111001010001111010111000011;
//0.2
inputlayer[5][0][0]=32'b00111110010011001100110011001101;
//0.2
inputlayer[6][0][0]=32'b00111110100110011001100110011010;
//0.7
inputlayer[7][0][0]=32'b00111111001100110011001100110011;
//-0.2
inputlayer[8][0][0]=32'b10111110010011001100110011001101;
//1
inputlayer[9][0][0]=32'b00111111100000000000000000000000;
#600
//-0.24
inputlayer[0][0][0]=32'b10111110011101011100001010001111;
//1
inputlayer[1][0][0]=32'b00111111100000000000000000000000;
//-1
inputlayer[2][0][0]=32'b10111111100000000000000000000000;
//0.5
inputlayer[3][0][0]=32'b00111111000000000000000000000000;
//-0.5
inputlayer[4][0][0]=32'b10111111000000000000000000000000;
//0.2
inputlayer[5][0][0]=32'b00111110010011001100110011001101;
//-0.5
inputlayer[6][0][0]=32'b10111111000000000000000000000000;
//1
inputlayer[7][0][0]=32'b00111111100000000000000000000000;
//0
inputlayer[8][0][0]=32'b00000000000000000000000000000000;
//0.3
inputlayer[9][0][0]=32'b00111110100110011001100110011010;
#600
//-1
inputlayer[0][0][0]=32'b10111111100000000000000000000000;
//0.7
inputlayer[1][0][0]=32'b00111111001100110011001100110011;
//-0.5
inputlayer[2][0][0]=32'b10111111000000000000000000000000;
//0.5
inputlayer[3][0][0]=32'b00111111000000000000000000000000;
//-0.66
inputlayer[4][0][0]=32'b10111111001010001111010111000011;
//0.2
inputlayer[5][0][0]=32'b00111110010011001100110011001101;
//2
inputlayer[6][0][0]=32'b01000000000000000000000000000000;
//-1
inputlayer[7][0][0]=32'b10111111100000000000000000000000;
//-0.2
inputlayer[8][0][0]=32'b10111110010011001100110011001101;
//0.5
inputlayer[9][0][0]=32'b00111111000000000000000000000000;
#2400
$finish;
end
always begin
forever #300 clock = ~clock;
end
always@(negedge clock)
begin
#600;
end
endmodule