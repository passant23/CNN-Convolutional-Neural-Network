`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/07/2020 03:11:01 PM
// Design Name: 
// Module Name: avg_3D_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

include "avg_3D.sv";
module avg_3D_tb;
localparam Period = 0.1; 
reg [31:0] ImagesIn [3] [10][10]; 
reg     clk ,start;
wire [31:0] ImagesOut [3][5][5]; 
wire [31:0] tempImage [3][10][10];
// -------------- Image 1 ----------------------

assign tempImage [0][0][0]=32'b00111111100000000000000000000000;  assign tempImage[0][0][1]=32'b01000000000000000000000000000000; assign tempImage[0][0][2]=32'b01000000010000000000000000000000;  assign tempImage[0][0][3]=32'b01000000100000000000000000000000;
assign tempImage[0][0][4]=32'b01000000101000000000000000000000;  assign tempImage[0][0][5]=32'b01000000110000000000000000000000; assign tempImage[0][0][6]=32'b01000000111000000000000000000000;  assign tempImage[0][0][7]=32'b01000001000000000000000000000000;
assign tempImage[0][0][8]=32'b01000001000100000000000000000000;  assign tempImage[0][0][9]=32'b01000001001000000000000000000000; assign tempImage[0][1][0]=32'b01000001001100000000000000000000;  assign tempImage[0][1][1]=32'b01000001010000000000000000000000;
assign tempImage [0][1][2]=32'b01000001010100000000000000000000; assign tempImage[0][1][3]=32'b01000001011000000000000000000000; assign tempImage [0][1][4]=32'b01000001011100000000000000000000; assign tempImage[0][1][5]=32'b01000001100000000000000000000000;
assign tempImage[0][1][6]=32'b01000001100010000000000000000000;  assign tempImage[0][1][7]=32'b01000001100100000000000000000000; assign tempImage[0][1][8]=32'b01000001100110000000000000000000;  assign tempImage[0][1][9]=32'b01000001101000000000000000000000;
assign tempImage[0][2][0]=32'b01000001101010000000000000000000;  assign tempImage[0][2][1]=32'b01000001101100000000000000000000; assign tempImage[0][2][2]=32'b01000001101110000000000000000000;  assign tempImage[0][2][3]=32'b01000001110000000000000000000000;
assign tempImage[0][2][4]=32'b01000001110010000000000000000000;  
//
assign tempImage[0][2][5]=32'b00111111100000000000000000000000;  assign tempImage[0][2][6]=32'b01000000000000000000000000000000; assign tempImage[0][2][7]=32'b01000000010000000000000000000000;  assign tempImage[0][2][8]=32'b01000000100000000000000000000000;
assign tempImage[0][2][9]=32'b01000000101000000000000000000000;  assign tempImage[0][3][0]=32'b01000000110000000000000000000000; assign tempImage[0][3][1]=32'b01000000111000000000000000000000;  assign tempImage[0][3][2]=32'b01000001000000000000000000000000;
assign tempImage[0][3][3]=32'b01000001000100000000000000000000;  assign tempImage[0][3][4]=32'b01000001001000000000000000000000; assign tempImage[0][3][5]=32'b01000001001100000000000000000000;  assign tempImage[0][3][6]=32'b01000001010000000000000000000000;
assign tempImage[0] [3][7]=32'b01000001010100000000000000000000; assign tempImage[0][3][8]=32'b01000001011000000000000000000000; assign tempImage[0] [3][9]=32'b01000001011100000000000000000000; assign tempImage[0][4][0]=32'b01000001100000000000000000000000;
assign tempImage[0][4][1]=32'b01000001100010000000000000000000;  assign tempImage[0][4][2]=32'b01000001100100000000000000000000; assign tempImage[0][4][3]=32'b01000001100110000000000000000000;  assign tempImage[0] [4][4]=32'b01000001101000000000000000000000;
assign tempImage[0][4][5]=32'b01000001101010000000000000000000;  assign tempImage[0][4][6]=32'b01000001101100000000000000000000; assign tempImage[0][4][7]=32'b01000001101110000000000000000000;  assign tempImage[0][4][8]=32'b01000001110000000000000000000000;
assign tempImage[0][4][9]=32'b01000001110010000000000000000000;
//
assign tempImage[0][5][0]=32'b00111111100000000000000000000000;  assign tempImage[0][5][1]=32'b01000000000000000000000000000000; assign tempImage[0][5][2]=32'b01000000010000000000000000000000;  assign tempImage[0][5][3]=32'b01000000100000000000000000000000;
assign tempImage[0][5][4]=32'b01000000101000000000000000000000;  assign tempImage[0][5][5]=32'b01000000110000000000000000000000; assign tempImage[0][5][6]=32'b01000000111000000000000000000000;  assign tempImage[0][5][7]=32'b01000001000000000000000000000000;
assign tempImage[0][5][8]=32'b01000001000100000000000000000000;  assign tempImage[0][5][9]=32'b01000001001000000000000000000000; assign tempImage[0][6][0]=32'b01000001001100000000000000000000;  assign tempImage[0][6][1]=32'b01000001010000000000000000000000;
assign tempImage [0][6][2]=32'b01000001010100000000000000000000; assign tempImage[0][6][3]=32'b01000001011000000000000000000000; assign tempImage[0] [6][4]=32'b01000001011100000000000000000000; assign tempImage[0][6][5]=32'b01000001100000000000000000000000;
assign tempImage[0][6][6]=32'b01000001100010000000000000000000;  assign tempImage[0][6][7]=32'b01000001100100000000000000000000; assign tempImage[0][6][8]=32'b01000001100110000000000000000000;  assign tempImage[0][6][9]=32'b01000001101000000000000000000000;
assign tempImage[0][7][0]=32'b01000001101010000000000000000000;  assign tempImage[0][7][1]=32'b01000001101100000000000000000000; assign tempImage[0][7][2]=32'b01000001101110000000000000000000;  assign tempImage[0][7][3]=32'b01000001110000000000000000000000;
assign tempImage[0][7][4]=32'b01000001110010000000000000000000;  
//
assign tempImage[0][7][5]=32'b00111111100000000000000000000000;  assign tempImage[0][7][6]=32'b01000000000000000000000000000000; assign tempImage[0][7][7]=32'b01000000010000000000000000000000;  assign tempImage[0][7][8]=32'b01000000100000000000000000000000;
assign tempImage[0][7][9]=32'b01000000101000000000000000000000;  assign tempImage[0][8][0]=32'b01000000110000000000000000000000; assign tempImage[0][8][1]=32'b01000000111000000000000000000000;  assign tempImage[0][8][2]=32'b01000001000000000000000000000000;
assign tempImage[0][8][3]=32'b01000001000100000000000000000000;  assign tempImage[0][8][4]=32'b01000001001000000000000000000000; assign tempImage[0][8][5]=32'b01000001001100000000000000000000;  assign tempImage[0][8][6]=32'b01000001010000000000000000000000;
assign tempImage[0][8][7]=32'b01000001010100000000000000000000;  assign tempImage[0][8][8]=32'b01000001011000000000000000000000; assign tempImage[0] [8][9]=32'b01000001011100000000000000000000; assign tempImage[0][9][0]=32'b01000001100000000000000000000000;
assign tempImage[0][9][1]=32'b01000001100010000000000000000000;  assign tempImage[0][9][2]=32'b01000001100100000000000000000000; assign tempImage[0][9][3]=32'b01000001100110000000000000000000;  assign tempImage[0][9][4]=32'b01000001101000000000000000000000;
assign tempImage[0][9][5]=32'b01000001101010000000000000000000;  assign tempImage[0][9][6]=32'b01000001101100000000000000000000; assign tempImage[0][9][7]=32'b01000001101110000000000000000000;  assign tempImage[0][9][8]=32'b01000001110000000000000000000000;
assign tempImage[0][9][9]=32'b01000001110010000000000000000000;

// -------------- Image 2 ----------------------

assign tempImage [1][0][0]=32'b00111111100000000000000000000000;  assign tempImage[1][0][1]=32'b01000000000000000000000000000000; assign tempImage[1][0][2]=32'b01000000010000000000000000000000;  assign tempImage[1][0][3]=32'b01000000100000000000000000000000;
assign tempImage[1][0][4]=32'b01000000101000000000000000000000;  assign tempImage[1][0][5]=32'b01000000110000000000000000000000; assign tempImage[1][0][6]=32'b01000000111000000000000000000000;  assign tempImage[1][0][7]=32'b01000001000000000000000000000000;
assign tempImage[1][0][8]=32'b01000001000100000000000000000000;  assign tempImage[1][0][9]=32'b01000001001000000000000000000000; assign tempImage[1][1][0]=32'b01000001001100000000000000000000;  assign tempImage[1][1][1]=32'b01000001010000000000000000000000;
assign tempImage [1][1][2]=32'b01000001010100000000000000000000; assign tempImage[1][1][3]=32'b01000001011000000000000000000000; assign tempImage [1][1][4]=32'b01000001011100000000000000000000; assign tempImage[1][1][5]=32'b01000001100000000000000000000000;
assign tempImage[1][1][6]=32'b01000001100010000000000000000000;  assign tempImage[1][1][7]=32'b01000001100100000000000000000000; assign tempImage[1][1][8]=32'b01000001100110000000000000000000;  assign tempImage[1][1][9]=32'b01000001101000000000000000000000;
assign tempImage[1][2][0]=32'b01000001101010000000000000000000;  assign tempImage[1][2][1]=32'b01000001101100000000000000000000; assign tempImage[1][2][2]=32'b01000001101110000000000000000000;  assign tempImage[1][2][3]=32'b01000001110000000000000000000000;
assign tempImage[1][2][4]=32'b01000001110010000000000000000000;  
//
assign tempImage[1][2][5]=32'b00111111100000000000000000000000;  assign tempImage[1][2][6]=32'b01000000000000000000000000000000; assign tempImage[1][2][7]=32'b01000000010000000000000000000000;  assign tempImage[1][2][8]=32'b01000000100000000000000000000000;
assign tempImage[1][2][9]=32'b01000000101000000000000000000000;  assign tempImage[1][3][0]=32'b01000000110000000000000000000000; assign tempImage[1][3][1]=32'b01000000111000000000000000000000;  assign tempImage[1][3][2]=32'b01000001000000000000000000000000;
assign tempImage[1][3][3]=32'b01000001000100000000000000000000;  assign tempImage[1][3][4]=32'b01000001001000000000000000000000; assign tempImage[1][3][5]=32'b01000001001100000000000000000000;  assign tempImage[1][3][6]=32'b01000001010000000000000000000000;
assign tempImage[1] [3][7]=32'b01000001010100000000000000000000; assign tempImage[1][3][8]=32'b01000001011000000000000000000000; assign tempImage[1] [3][9]=32'b01000001011100000000000000000000; assign tempImage[1][4][0]=32'b01000001100000000000000000000000;
assign tempImage[1][4][1]=32'b01000001100010000000000000000000;  assign tempImage[1][4][2]=32'b01000001100100000000000000000000; assign tempImage[1][4][3]=32'b01000001100110000000000000000000;  assign tempImage[1] [4][4]=32'b01000001101000000000000000000000;
assign tempImage[1][4][5]=32'b01000001101010000000000000000000;  assign tempImage[1][4][6]=32'b01000001101100000000000000000000; assign tempImage[1][4][7]=32'b01000001101110000000000000000000;  assign tempImage[1][4][8]=32'b01000001110000000000000000000000;
assign tempImage[1][4][9]=32'b01000001110010000000000000000000;
//
assign tempImage[1][5][0]=32'b00111111100000000000000000000000;  assign tempImage[1][5][1]=32'b01000000000000000000000000000000; assign tempImage[1][5][2]=32'b01000000010000000000000000000000;  assign tempImage[1][5][3]=32'b01000000100000000000000000000000;
assign tempImage[1][5][4]=32'b01000000101000000000000000000000;  assign tempImage[1][5][5]=32'b01000000110000000000000000000000; assign tempImage[1][5][6]=32'b01000000111000000000000000000000;  assign tempImage[1][5][7]=32'b01000001000000000000000000000000;
assign tempImage[1][5][8]=32'b01000001000100000000000000000000;  assign tempImage[1][5][9]=32'b01000001001000000000000000000000; assign tempImage[1][6][0]=32'b01000001001100000000000000000000;  assign tempImage[1][6][1]=32'b01000001010000000000000000000000;
assign tempImage [1][6][2]=32'b01000001010100000000000000000000; assign tempImage[1][6][3]=32'b01000001011000000000000000000000; assign tempImage[1] [6][4]=32'b01000001011100000000000000000000; assign tempImage[1][6][5]=32'b01000001100000000000000000000000;
assign tempImage[1][6][6]=32'b01000001100010000000000000000000;  assign tempImage[1][6][7]=32'b01000001100100000000000000000000; assign tempImage[1][6][8]=32'b01000001100110000000000000000000;  assign tempImage[1][6][9]=32'b01000001101000000000000000000000;
assign tempImage[1][7][0]=32'b01000001101010000000000000000000;  assign tempImage[1][7][1]=32'b01000001101100000000000000000000; assign tempImage[1][7][2]=32'b01000001101110000000000000000000;  assign tempImage[1][7][3]=32'b01000001110000000000000000000000;
assign tempImage[1][7][4]=32'b01000001110010000000000000000000;  
//
assign tempImage[1][7][5]=32'b00111111100000000000000000000000;  assign tempImage[1][7][6]=32'b01000000000000000000000000000000; assign tempImage[1][7][7]=32'b01000000010000000000000000000000;  assign tempImage[1][7][8]=32'b01000000100000000000000000000000;
assign tempImage[1][7][9]=32'b01000000101000000000000000000000;  assign tempImage[1][8][0]=32'b01000000110000000000000000000000; assign tempImage[1][8][1]=32'b01000000111000000000000000000000;  assign tempImage[1][8][2]=32'b01000001000000000000000000000000;
assign tempImage[1][8][3]=32'b01000001000100000000000000000000;  assign tempImage[1][8][4]=32'b01000001001000000000000000000000; assign tempImage[1][8][5]=32'b01000001001100000000000000000000;  assign tempImage[1][8][6]=32'b01000001010000000000000000000000;
assign tempImage[1][8][7]=32'b01000001010100000000000000000000;  assign tempImage[1][8][8]=32'b01000001011000000000000000000000; assign tempImage[1] [8][9]=32'b01000001011100000000000000000000; assign tempImage[1][9][0]=32'b01000001100000000000000000000000;
assign tempImage[1][9][1]=32'b01000001100010000000000000000000;  assign tempImage[1][9][2]=32'b01000001100100000000000000000000; assign tempImage[1][9][3]=32'b01000001100110000000000000000000;  assign tempImage[1][9][4]=32'b01000001101000000000000000000000;
assign tempImage[1][9][5]=32'b01000001101010000000000000000000;  assign tempImage[1][9][6]=32'b01000001101100000000000000000000; assign tempImage[1][9][7]=32'b01000001101110000000000000000000;  assign tempImage[1][9][8]=32'b01000001110000000000000000000000;
assign tempImage[1][9][9]=32'b01000001110010000000000000000000;

// -------------- Image 3 ----------------------
assign tempImage [2][0][0]=32'b00111111100000000000000000000000;  assign tempImage[2][0][1]=32'b01000000000000000000000000000000; assign tempImage[2][0][2]=32'b01000000010000000000000000000000;  assign tempImage[2][0][3]=32'b01000000100000000000000000000000;
assign tempImage[2][0][4]=32'b01000000101000000000000000000000;  assign tempImage[2][0][5]=32'b01000000110000000000000000000000; assign tempImage[2][0][6]=32'b01000000111000000000000000000000;  assign tempImage[2][0][7]=32'b01000001000000000000000000000000;
assign tempImage[2][0][8]=32'b01000001000100000000000000000000;  assign tempImage[2][0][9]=32'b01000001001000000000000000000000; assign tempImage[2][1][0]=32'b01000001001100000000000000000000;  assign tempImage[2][1][1]=32'b01000001010000000000000000000000;
assign tempImage [2][1][2]=32'b01000001010100000000000000000000; assign tempImage[2][1][3]=32'b01000001011000000000000000000000; assign tempImage [2][1][4]=32'b01000001011100000000000000000000; assign tempImage[2][1][5]=32'b01000001100000000000000000000000;
assign tempImage[2][1][6]=32'b01000001100010000000000000000000;  assign tempImage[2][1][7]=32'b01000001100100000000000000000000; assign tempImage[2][1][8]=32'b01000001100110000000000000000000;  assign tempImage[2][1][9]=32'b01000001101000000000000000000000;
assign tempImage[2][2][0]=32'b01000001101010000000000000000000;  assign tempImage[2][2][1]=32'b01000001101100000000000000000000; assign tempImage[2][2][2]=32'b01000001101110000000000000000000;  assign tempImage[2][2][3]=32'b01000001110000000000000000000000;
assign tempImage[2][2][4]=32'b01000001110010000000000000000000;  
//
assign tempImage[2][2][5]=32'b00111111100000000000000000000000;  assign tempImage[2][2][6]=32'b01000000000000000000000000000000; assign tempImage[2][2][7]=32'b01000000010000000000000000000000;  assign tempImage[2][2][8]=32'b01000000100000000000000000000000;
assign tempImage[2][2][9]=32'b01000000101000000000000000000000;  assign tempImage[2][3][0]=32'b01000000110000000000000000000000; assign tempImage[2][3][1]=32'b01000000111000000000000000000000;  assign tempImage[2][3][2]=32'b01000001000000000000000000000000;
assign tempImage[2][3][3]=32'b01000001000100000000000000000000;  assign tempImage[2][3][4]=32'b01000001001000000000000000000000; assign tempImage[2][3][5]=32'b01000001001100000000000000000000;  assign tempImage[2][3][6]=32'b01000001010000000000000000000000;
assign tempImage[2] [3][7]=32'b01000001010100000000000000000000; assign tempImage[2][3][8]=32'b01000001011000000000000000000000; assign tempImage[2] [3][9]=32'b01000001011100000000000000000000; assign tempImage[2][4][0]=32'b01000001100000000000000000000000;
assign tempImage[2][4][1]=32'b01000001100010000000000000000000;  assign tempImage[2][4][2]=32'b01000001100100000000000000000000; assign tempImage[2][4][3]=32'b01000001100110000000000000000000;  assign tempImage[2] [4][4]=32'b01000001101000000000000000000000;
assign tempImage[2][4][5]=32'b01000001101010000000000000000000;  assign tempImage[2][4][6]=32'b01000001101100000000000000000000; assign tempImage[2][4][7]=32'b01000001101110000000000000000000;  assign tempImage[2][4][8]=32'b01000001110000000000000000000000;
assign tempImage[2][4][9]=32'b01000001110010000000000000000000;
//
assign tempImage[2][5][0]=32'b00111111100000000000000000000000;  assign tempImage[2][5][1]=32'b01000000000000000000000000000000; assign tempImage[2][5][2]=32'b01000000010000000000000000000000;  assign tempImage[2][5][3]=32'b01000000100000000000000000000000;
assign tempImage[2][5][4]=32'b01000000101000000000000000000000;  assign tempImage[2][5][5]=32'b01000000110000000000000000000000; assign tempImage[2][5][6]=32'b01000000111000000000000000000000;  assign tempImage[2][5][7]=32'b01000001000000000000000000000000;
assign tempImage[2][5][8]=32'b01000001000100000000000000000000;  assign tempImage[2][5][9]=32'b01000001001000000000000000000000; assign tempImage[2][6][0]=32'b01000001001100000000000000000000;  assign tempImage[2][6][1]=32'b01000001010000000000000000000000;
assign tempImage [2][6][2]=32'b01000001010100000000000000000000; assign tempImage[2][6][3]=32'b01000001011000000000000000000000; assign tempImage[2] [6][4]=32'b01000001011100000000000000000000; assign tempImage[2][6][5]=32'b01000001100000000000000000000000;
assign tempImage[2][6][6]=32'b01000001100010000000000000000000;  assign tempImage[2][6][7]=32'b01000001100100000000000000000000; assign tempImage[2][6][8]=32'b01000001100110000000000000000000;  assign tempImage[2][6][9]=32'b01000001101000000000000000000000;
assign tempImage[2][7][0]=32'b01000001101010000000000000000000;  assign tempImage[2][7][1]=32'b01000001101100000000000000000000; assign tempImage[2][7][2]=32'b01000001101110000000000000000000;  assign tempImage[2][7][3]=32'b01000001110000000000000000000000;
assign tempImage[2][7][4]=32'b01000001110010000000000000000000;  
//
assign tempImage[2][7][5]=32'b00111111100000000000000000000000;  assign tempImage[2][7][6]=32'b01000000000000000000000000000000; assign tempImage[2][7][7]=32'b01000000010000000000000000000000;  assign tempImage[2][7][8]=32'b01000000100000000000000000000000;
assign tempImage[2][7][9]=32'b01000000101000000000000000000000;  assign tempImage[2][8][0]=32'b01000000110000000000000000000000; assign tempImage[2][8][1]=32'b01000000111000000000000000000000;  assign tempImage[2][8][2]=32'b01000001000000000000000000000000;
assign tempImage[2][8][3]=32'b01000001000100000000000000000000;  assign tempImage[2][8][4]=32'b01000001001000000000000000000000; assign tempImage[2][8][5]=32'b01000001001100000000000000000000;  assign tempImage[2][8][6]=32'b01000001010000000000000000000000;
assign tempImage[2][8][7]=32'b01000001010100000000000000000000;  assign tempImage[2][8][8]=32'b01000001011000000000000000000000; assign tempImage[2] [8][9]=32'b01000001011100000000000000000000; assign tempImage[2][9][0]=32'b01000001100000000000000000000000;
assign tempImage[2][9][1]=32'b01000001100010000000000000000000;  assign tempImage[2][9][2]=32'b01000001100100000000000000000000; assign tempImage[2][9][3]=32'b01000001100110000000000000000000;  assign tempImage[2][9][4]=32'b01000001101000000000000000000000;
assign tempImage[2][9][5]=32'b01000001101010000000000000000000;  assign tempImage[2][9][6]=32'b01000001101100000000000000000000; assign tempImage[2][9][7]=32'b01000001101110000000000000000000;  assign tempImage[2][9][8]=32'b01000001110000000000000000000000;
assign tempImage[2][9][9]=32'b01000001110010000000000000000000;
// -------------------------------------------------------------------- //

 always
    begin
    #(Period/2) clk = ~clk;
    end
initial
  begin
   start=0;
   clk=0;
   //#(Period/2) //  1st Rising edge: Assign pixel of image
   ImagesIn=tempImage; 
   #Period // Next Falling edge
   start=1;
   #(126*Period)
   $stop;
   end
      
avg_3D images (
.ImagesIn(ImagesIn),
.clk(clk),
.start(start),
.ImagesOut(ImagesOut)
);
endmodule
