`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/09/2020 09:07:07 PM
// Design Name: 
// Module Name: testbench_SoftmaxMaxIndex
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module testbench_SoftmaxMaxIndex();
 parameter datawidth=32;
   reg clock;
   reg reset;
   reg [datawidth-1:0] inputS [10][1][1];  
   wire [datawidth-1:0] outputS [10][1][1];
   wire [datawidth-1:0] max_S;
   wire [3:0] index_S;
   wire done;
   
 softmax_max_index softmax_integrated (clock,reset,inputS,outputS,max_S,index_S,done);
   
   
   initial begin
   clock=1'b1;
   reset=1'b0;
   //0
   inputS[0][0][0]=32'b00000000000000000000000000000000;
   //1
   inputS[1][0][0]=32'b00111111100000000000000000000000;
   //-1
   inputS[2][0][0]=32'b10111111100000000000000000000000;
   //0.5
   inputS[3][0][0]=32'b00111111000000000000000000000000;
   //1
   inputS[4][0][0]=32'b00111111100000000000000000000000;
   //0.2
   inputS[5][0][0]=32'b00111110010011001100110011001101;
   //-0.5
   inputS[6][0][0]=32'b10111111000000000000000000000000;
   //0.3
   inputS[7][0][0]=32'b00111110100110011001100110011010;
   //0
   inputS[8][0][0]=32'b00000000000000000000000000000000;
   //0.7
   inputS[9][0][0]=32'b00111111001100110011001100110011;
   #600
   //-1
   inputS[0][0][0]=32'b10111111100000000000000000000000;
   //0
   inputS[1][0][0]=32'b00000000000000000000000000000000;
   //-0.5
   inputS[2][0][0]=32'b10111111000000000000000000000000;
   //0.5
   inputS[3][0][0]=32'b00111111000000000000000000000000;
   //-0.66
   inputS[4][0][0]=32'b10111111001010001111010111000011;
   //0.2
   inputS[5][0][0]=32'b00111110010011001100110011001101;
   //0.2
   inputS[6][0][0]=32'b00111110100110011001100110011010;
   //0.7
   inputS[7][0][0]=32'b00111111001100110011001100110011;
   //-0.2
   inputS[8][0][0]=32'b10111110010011001100110011001101;
   //1
   inputS[9][0][0]=32'b00111111100000000000000000000000;
   #600
   //-0.24
   inputS[0][0][0]=32'b10111110011101011100001010001111;
   //1
   inputS[1][0][0]=32'b00111111100000000000000000000000;
   //-1
   inputS[2][0][0]=32'b10111111100000000000000000000000;
   //0.5
   inputS[3][0][0]=32'b00111111000000000000000000000000;
   //-0.5
   inputS[4][0][0]=32'b10111111000000000000000000000000;
   //0.2
   inputS[5][0][0]=32'b00111110010011001100110011001101;
   //-0.5
   inputS[6][0][0]=32'b10111111000000000000000000000000;
   //1
   inputS[7][0][0]=32'b00111111100000000000000000000000;
   //0
   inputS[8][0][0]=32'b00000000000000000000000000000000;
   //0.3
   inputS[9][0][0]=32'b00111110100110011001100110011010;
   #600
   //-1
   inputS[0][0][0]=32'b10111111100000000000000000000000;
   //0.7
   inputS[1][0][0]=32'b00111111001100110011001100110011;
   //-0.5
   inputS[2][0][0]=32'b10111111000000000000000000000000;
   //0.5
   inputS[3][0][0]=32'b00111111000000000000000000000000;
   //-0.66
   inputS[4][0][0]=32'b10111111001010001111010111000011;
   //0.2
   inputS[5][0][0]=32'b00111110010011001100110011001101;
   //2
   inputS[6][0][0]=32'b01000000000000000000000000000000;
   //-1
   inputS[7][0][0]=32'b10111111100000000000000000000000;
   //-0.2
   inputS[8][0][0]=32'b10111110010011001100110011001101;
   //0.5
   inputS[9][0][0]=32'b00111111000000000000000000000000;
   #2400
   $finish;
   end
   always begin
   forever #300 clock = ~clock;
   end
   always@(negedge clock)
   begin
   #600;
   end

endmodule