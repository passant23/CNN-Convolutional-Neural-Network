`timescale 1ns / 1ps
module testbench_comparingSoftmax();
parameter datawidth=32;
reg clock;
reg [datawidth-1:0] softmax_out [9:0][1][1];  
wire [datawidth-1:0] max_out;
wire [3:0] max_index;

comparingSoftmax cm(clock,softmax_out,max_out,max_index);
initial begin
clock=1'b1;
//e^1
softmax_out[0][0][0]=32'b01000000001011010111000010100100;
//e^0
softmax_out[1][0][0]=32'b00111111100000000000000000000000;
//e^-0.5
softmax_out[2][0][0]=32'b00111111000110110100001110010110;
//e^0.5
softmax_out[3][0][0]=32'b00111111110100110000100010011010;
//e^0
softmax_out[4][0][0]=32'b00111111010100011001011001010011;
//e^-0.2
softmax_out[5][0][0]=32'b00111111010100011001011001010011;
//e^0.4
softmax_out[6][0][0]=32'b00111111101111101111001101001101;
//e^-1
softmax_out[7][0][0]=32'b00111110101111000101000001001000;
//e^0.7
softmax_out[8][0][0]=32'b01000000000000001110000001110110;
//e^0.9
softmax_out[9][0][0]=32'b01000000000111010110101000010110;
#30
//e^-1
softmax_out[0][0][0]=32'b00111110101111000101000001001000;
//e^0
softmax_out[1][0][0]=32'b00111111100000000000000000000000;
//e^-1
softmax_out[2][0][0]=32'b00111110101111000101000001001000;
//e^0.5
softmax_out[3][0][0]=32'b00111111110100110000100010011010;
//e^0.7
softmax_out[4][0][0]=32'b01000000000000001110000001110110;
//e^-0.2
softmax_out[5][0][0]=32'b00111111010100011001011001010011;
//e^-0.5
softmax_out[6][0][0]=32'b00111111000110110100001110010110;
//e^0.9
softmax_out[7][0][0]=32'b01000000000111010110101000010110;
//e^0.7
softmax_out[8][0][0]=32'b01000000000000001110000001110110;
//e^-0.2
softmax_out[9][0][0]=32'b00111111010100011001011001010011;
#30
//e^-0.5
softmax_out[0][0][0]=32'b00111111000110110100001110010110;
//e^0
softmax_out[1][0][0]=32'b00111111100000000000000000000000;
//e^1
softmax_out[2][0][0]=32'b01000000001011010111000010100100;
//e^0.6
softmax_out[3][0][0]=32'b00111111111010010011011101001100;
//e^0.3
softmax_out[4][0][0]=32'b00111111101011001100011000111111;
//e^-0.2
softmax_out[5][0][0]=32'b00111111010100011001011001010011;
//e^0.4
softmax_out[6][0][0]=32'b00111111101111101111001101001101;
//e^-1
softmax_out[7][0][0]=32'b00111110101111000101000001001000;
//e^0.7
softmax_out[8][0][0]=32'b01000000000000001110000001110110;
//e^0.9
softmax_out[9][0][0]=32'b01000000000111010110101000010110;
#120
$finish;
end
always begin
forever #15 clock = ~clock;
end
always@(negedge clock)
begin
#30;
end
endmodule