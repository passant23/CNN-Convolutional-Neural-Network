`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/30/2020 10:08:17 PM
// Design Name: 
// Module Name: avg_2D_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

include "AvgLayer.sv";
module avg_2D_tb;
// Setting the clock //
localparam Period = 0.1; 
reg [31:0] Imagein [10][10];
reg clk,start;
reg [31:0] tempImage [10][10];
wire [31:0] Imageout [5][5];
assign tempImage[0][0]=32'b00111111100000000000000000000000;  assign tempImage[0][1]=32'b01000000000000000000000000000000; assign tempImage[0][2]=32'b01000000010000000000000000000000;  assign tempImage[0][3]=32'b01000000100000000000000000000000;
assign tempImage[0][4]=32'b01000000101000000000000000000000;  assign tempImage[0][5]=32'b01000000110000000000000000000000; assign tempImage[0][6]=32'b01000000111000000000000000000000;  assign tempImage[0][7]=32'b01000001000000000000000000000000;
assign tempImage[0][8]=32'b01000001000100000000000000000000;  assign tempImage[0][9]=32'b01000001001000000000000000000000; assign tempImage[1][0]=32'b01000001001100000000000000000000;  assign tempImage[1][1]=32'b01000001010000000000000000000000;
assign tempImage [1][2]=32'b01000001010100000000000000000000; assign tempImage[1][3]=32'b01000001011000000000000000000000; assign tempImage [1][4]=32'b01000001011100000000000000000000; assign tempImage[1][5]=32'b01000001100000000000000000000000;
assign tempImage[1][6]=32'b01000001100010000000000000000000;  assign tempImage[1][7]=32'b01000001100100000000000000000000; assign tempImage[1][8]=32'b01000001100110000000000000000000;  assign tempImage[1][9]=32'b01000001101000000000000000000000;
assign tempImage[2][0]=32'b01000001101010000000000000000000;  assign tempImage[2][1]=32'b01000001101100000000000000000000; assign tempImage[2][2]=32'b01000001101110000000000000000000;  assign tempImage[2][3]=32'b01000001110000000000000000000000;
assign tempImage[2][4]=32'b01000001110010000000000000000000;  
//
assign tempImage[2][5]=32'b00111111100000000000000000000000;  assign tempImage[2][6]=32'b01000000000000000000000000000000; assign tempImage[2][7]=32'b01000000010000000000000000000000;  assign tempImage[2][8]=32'b01000000100000000000000000000000;
assign tempImage[2][9]=32'b01000000101000000000000000000000;  assign tempImage[3][0]=32'b01000000110000000000000000000000; assign tempImage[3][1]=32'b01000000111000000000000000000000;  assign tempImage[3][2]=32'b01000001000000000000000000000000;
assign tempImage[3][3]=32'b01000001000100000000000000000000;  assign tempImage[3][4]=32'b01000001001000000000000000000000; assign tempImage[3][5]=32'b01000001001100000000000000000000;  assign tempImage[3][6]=32'b01000001010000000000000000000000;
assign tempImage [3][7]=32'b01000001010100000000000000000000; assign tempImage[3][8]=32'b01000001011000000000000000000000; assign tempImage [3][9]=32'b01000001011100000000000000000000; assign tempImage[4][0]=32'b01000001100000000000000000000000;
assign tempImage[4][1]=32'b01000001100010000000000000000000;  assign tempImage[4][2]=32'b01000001100100000000000000000000; assign tempImage[4][3]=32'b01000001100110000000000000000000;  assign tempImage[4][4]=32'b01000001101000000000000000000000;
assign tempImage[4][5]=32'b01000001101010000000000000000000;  assign tempImage[4][6]=32'b01000001101100000000000000000000; assign tempImage[4][7]=32'b01000001101110000000000000000000;  assign tempImage[4][8]=32'b01000001110000000000000000000000;
assign tempImage[4][9]=32'b01000001110010000000000000000000;
//
assign tempImage[5][0]=32'b00111111100000000000000000000000;  assign tempImage[5][1]=32'b01000000000000000000000000000000; assign tempImage[5][2]=32'b01000000010000000000000000000000;  assign tempImage[5][3]=32'b01000000100000000000000000000000;
assign tempImage[5][4]=32'b01000000101000000000000000000000;  assign tempImage[5][5]=32'b01000000110000000000000000000000; assign tempImage[5][6]=32'b01000000111000000000000000000000;  assign tempImage[5][7]=32'b01000001000000000000000000000000;
assign tempImage[5][8]=32'b01000001000100000000000000000000;  assign tempImage[5][9]=32'b01000001001000000000000000000000; assign tempImage[6][0]=32'b01000001001100000000000000000000;  assign tempImage[6][1]=32'b01000001010000000000000000000000;
assign tempImage [6][2]=32'b01000001010100000000000000000000; assign tempImage[6][3]=32'b01000001011000000000000000000000; assign tempImage [6][4]=32'b01000001011100000000000000000000; assign tempImage[6][5]=32'b01000001100000000000000000000000;
assign tempImage[6][6]=32'b01000001100010000000000000000000;  assign tempImage[6][7]=32'b01000001100100000000000000000000; assign tempImage[6][8]=32'b01000001100110000000000000000000;  assign tempImage[6][9]=32'b01000001101000000000000000000000;
assign tempImage[7][0]=32'b01000001101010000000000000000000;  assign tempImage[7][1]=32'b01000001101100000000000000000000; assign tempImage[7][2]=32'b01000001101110000000000000000000;  assign tempImage[7][3]=32'b01000001110000000000000000000000;
assign tempImage[7][4]=32'b01000001110010000000000000000000;  
//
assign tempImage[7][5]=32'b00111111100000000000000000000000;  assign tempImage[7][6]=32'b01000000000000000000000000000000; assign tempImage[7][7]=32'b01000000010000000000000000000000;  assign tempImage[7][8]=32'b01000000100000000000000000000000;
assign tempImage[7][9]=32'b01000000101000000000000000000000;  assign tempImage[8][0]=32'b01000000110000000000000000000000; assign tempImage[8][1]=32'b01000000111000000000000000000000;  assign tempImage[8][2]=32'b01000001000000000000000000000000;
assign tempImage[8][3]=32'b01000001000100000000000000000000;  assign tempImage[8][4]=32'b01000001001000000000000000000000; assign tempImage[8][5]=32'b01000001001100000000000000000000;  assign tempImage[8][6]=32'b01000001010000000000000000000000;
assign tempImage [8][7]=32'b01000001010100000000000000000000; assign tempImage[8][8]=32'b01000001011000000000000000000000; assign tempImage [8][9]=32'b01000001011100000000000000000000; assign tempImage[9][0]=32'b01000001100000000000000000000000;
assign tempImage[9][1]=32'b01000001100010000000000000000000;  assign tempImage[9][2]=32'b01000001100100000000000000000000; assign tempImage[9][3]=32'b01000001100110000000000000000000;  assign tempImage[9][4]=32'b01000001101000000000000000000000;
assign tempImage[9][5]=32'b01000001101010000000000000000000;  assign tempImage[9][6]=32'b01000001101100000000000000000000; assign tempImage[9][7]=32'b01000001101110000000000000000000;  assign tempImage[9][8]=32'b01000001110000000000000000000000;
assign tempImage[9][9]=32'b01000001110010000000000000000000;
//

AvgLayer avg(
.ImageIn(Imagein),
.ImageOut(Imageout),
.start(start),
.clk(clk)
);
      always
      begin
      #(Period/2) clk = ~clk;
      end
initial
begin
start=0;
clk=0;
//#(Period/2) //  1st Rising edge: Assign pixel of image
Imagein=tempImage; 
#Period // Next Falling edge
start=1;
#(126*Period)
$stop;
end

endmodule

